module or3(input a,input b,input c,output y);
	or(y,a,b,c);
endmodule
