module not_gate(input a, output y);
    not(y, a);
endmodule
