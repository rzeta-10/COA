module xnor_gate(input a,input b,output y);
    xnor(y,a,b);
endmodule