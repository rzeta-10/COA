// and3.v
module and3(input a, input b, input c, output y);
    and(y, a, b, c);
endmodule