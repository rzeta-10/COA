module nor_gate(input a,input b,output y);
    nor(y,a,b);
endmodule